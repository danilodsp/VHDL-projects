LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY pacemaker IS
	PORT(
	
	);
END pacemaker;
