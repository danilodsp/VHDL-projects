LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY controller IS
	PORT(
	clk: IN STD_LOGIC;
	
	);
END controller;

ARCHITECTURE c_mp OF controller IS



END c_mp;
